package my_pack;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "sequence_item.sv"
    `include "fixed_write_sequence.sv"
    `include "fixed_write_read_sequence.sv"
    `include "incr_write_sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "environment.sv"
    `include "fixed_write_test.sv"
    `include "fixed_write_read_test.sv"
    `include "incr_write_test.sv"
    

endpackage
